module MCP0832(clk_out,in,di,cs);



endmodule
