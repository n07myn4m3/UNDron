/* -----------------------------------------------------
   wb_everloop
   -----------------------------------------------------
	██╗   ██╗███╗   ██╗██████╗ ██████╗  ██████╗ ███╗   ██╗    
	██║   ██║████╗  ██║██╔══██╗██╔══██╗██╔═══██╗████╗  ██║    
	██║   ██║██╔██╗ ██║██║  ██║██████╔╝██║   ██║██╔██╗ ██║    
	██║   ██║██║╚██╗██║██║  ██║██╔══██╗██║   ██║██║╚██╗██║    
	╚██████╔╝██║ ╚████║██████╔╝██║  ██║╚██████╔╝██║ ╚████║    
	 ╚═════╝ ╚═╝  ╚═══╝╚═════╝ ╚═╝  ╚═╝ ╚═════╝ ╚═╝  ╚═══╝  
   DESCRIPCIÓN DE LOS REGISTROS
   0x00 everloop_ram

   FUNCIONAMIENTO
   * La direccion adr_a de la memoria RAM depende de la direccion escrita presente en el wishbone
     y de un valor de uno o cero 
   * ---   

   CONVENCIONES      
   * --- 
   * ---

   INDICADORES
   * PROBLEMA: Situacion que genera conflicto y debe corregirse
   * NPI: Declaracion que no se conoce
*/

module wb_everloop#(
  parameter mem_file_name = "none"  
)(
  input              clk,
  input              rst,
     
   // Wishbone interface
   input              wb_stb_i,
   input              wb_cyc_i,
   output             wb_ack_o,
   input              wb_we_i,
   input       [31:0] wb_adr_i,
   input        [3:0] wb_sel_i,
   input       [31:0] wb_dat_i,
   output reg  [31:0] wb_dat_o,

   // Everloop interface
   output everloop_led_ctl // Es la salida que va conectada al everloop fisico
   //input  led_fb,  // Esta entrada no es utilizada NPI
);


assign wb_ack_o = wb_stb_i & wb_cyc_i & ack;

wire wb_rd = wb_stb_i & wb_cyc_i & ~wb_we_i;
wire wb_wr = wb_stb_i & wb_cyc_i &  wb_we_i;
reg  ack;


// Al parecer son cables y registros usados por las memorias
wire [7:0]  data_b;
wire [10:0] adr_b;
reg  [2:0]  swr; // NPI
reg  [7:0]  data_a;
reg         add_adr_a; // NPI

always @(negedge clk)  swr <= {swr[1:0],wb_wr};

wire wr_fallingedge = (swr[2:1]==2'b10);



everloop everloop0(
  .clk(clk),
  .rst(rst),
  .address(adr_b),           // Se conecta a la memoria RAM de doble puerto 
  .data_RGB(data_b),
  .everloop_d(everloop_led_ctl)
);

everloop_ram #(
  .adr_width(11), 
  .dat_width(8), 
  .mem_file_name(mem_file_name)
) everloopram0(
  .clk_a(clk),
  .en_a (wb_wr | add_adr_a), // Solo habilita si el wishbone esta en modo de escritura y si el habilitador esta disponible
  .adr_a({wb_adr_i[9:0],add_adr_a}), 
  .dat_a(data_a[7:0]),
  .we_a (wb_wr | add_adr_a), // Solo escribe si el wishbone esta en modo de escritura y si el habilitador esta disponible
  .clk_b(clk),
  .en_b (1'b1),              //Por defecto se dejo habilitado la lectura de la memoria RAM
  .adr_b(adr_b),
  .dat_b(data_b)	
);

always @(posedge clk)
begin

case({wb_wr,wr_fallingedge}) //Solo si esta en modo de escritura y detecta un flanco de bajada
  2'b10: begin
    data_a    <= wb_dat_i;   //Un dato queda almacenado en data_a
    add_adr_a <= 0;          //No puedo escribirlo
  end
  2'b01:begin
    data_a    <= data_a >>8; //Desplazo el numero para que puedan observarse el siguiente byte
    add_adr_a <= 1;          //Envia la informacion a la memoria ram
  end
  
  default: begin
    data_a    <= data_a;
    add_adr_a <= 0;
  end
endcase
end

endmodule
